`default_nettype none
`include "def.sv"
module executer(
  input wire CLK,
  input control_info CTR_INFO,

  output
);


always @(posedge CLK) begin



end

end module
`default_nettype wire